magic
tech scmos
timestamp 1733078276
<< nwell >>
rect -30 -13 -6 21
rect 12 19 36 53
rect 45 18 79 42
rect 12 -66 36 -32
rect 104 -43 128 -9
<< ntransistor >>
rect 23 1 25 11
rect 115 1 117 11
rect -19 -31 -17 -21
rect 52 -50 62 -48
rect 23 -84 25 -74
<< ptransistor >>
rect 23 27 25 47
rect 53 29 73 31
rect -19 -5 -17 15
rect 115 -37 117 -17
rect 23 -58 25 -38
<< ndiffusion >>
rect 22 1 23 11
rect 25 1 26 11
rect 114 1 115 11
rect 117 1 118 11
rect -20 -31 -19 -21
rect -17 -31 -16 -21
rect 52 -48 62 -47
rect 52 -51 62 -50
rect 22 -84 23 -74
rect 25 -84 26 -74
<< pdiffusion >>
rect 22 27 23 47
rect 25 27 26 47
rect 53 31 73 32
rect 53 28 73 29
rect -20 -5 -19 15
rect -17 -5 -16 15
rect 114 -37 115 -17
rect 117 -37 118 -17
rect 22 -58 23 -38
rect 25 -58 26 -38
<< ndcontact >>
rect 18 1 22 11
rect 26 1 30 11
rect 110 1 114 11
rect 118 1 122 11
rect -24 -31 -20 -21
rect -16 -31 -12 -21
rect 52 -47 62 -43
rect 52 -55 62 -51
rect 18 -84 22 -74
rect 26 -84 30 -74
<< pdcontact >>
rect 18 27 22 47
rect 26 27 30 47
rect 53 32 73 36
rect -24 -5 -20 15
rect -16 -5 -12 15
rect 53 24 73 28
rect 110 -37 114 -17
rect 118 -37 122 -17
rect 18 -58 22 -38
rect 26 -58 30 -38
<< polysilicon >>
rect 23 47 25 50
rect 45 31 49 42
rect 45 29 53 31
rect 73 29 76 31
rect -19 15 -17 18
rect 23 11 25 27
rect 107 13 117 17
rect 115 11 117 13
rect 23 -2 25 1
rect 115 -2 117 1
rect -19 -21 -17 -5
rect 115 -14 122 -10
rect 115 -17 117 -14
rect -19 -34 -17 -31
rect 23 -38 25 -35
rect 115 -40 117 -37
rect 45 -50 52 -48
rect 62 -50 65 -48
rect 23 -74 25 -58
rect 23 -87 25 -84
<< polycontact >>
rect 45 42 49 46
rect 143 32 152 36
rect 19 14 23 18
rect 103 13 107 17
rect -23 -18 -19 -14
rect 122 -14 126 -10
rect 45 -54 49 -50
rect 19 -71 23 -67
<< metal1 >>
rect -43 52 49 56
rect -43 -14 -39 52
rect 18 47 22 52
rect 45 46 49 52
rect 47 24 53 28
rect -30 20 -6 24
rect -24 15 -20 20
rect 0 14 19 18
rect 0 -5 4 14
rect 47 -5 51 24
rect 102 1 110 5
rect 118 1 122 11
rect 0 -9 51 -5
rect -43 -18 -23 -14
rect -43 -89 -39 -18
rect 0 -26 4 -9
rect 0 -30 51 -26
rect -24 -36 -20 -31
rect -30 -40 -6 -36
rect 0 -67 4 -30
rect 47 -43 51 -30
rect 122 -37 129 -33
rect 47 -47 52 -43
rect 0 -71 19 -67
rect 18 -89 22 -84
rect 45 -89 49 -54
rect -43 -93 49 -89
<< metal2 >>
rect 26 18 30 47
rect 39 32 154 36
rect 39 18 43 32
rect -16 -14 -12 15
rect 26 14 43 18
rect 18 -14 22 11
rect 26 1 30 14
rect 79 13 107 17
rect -16 -18 22 -14
rect -16 -31 -12 -18
rect 18 -58 22 -18
rect 79 -33 83 13
rect 118 1 122 32
rect 131 -10 135 32
rect 122 -14 135 -10
rect 110 -33 114 -17
rect 79 -37 114 -33
rect 26 -67 30 -38
rect 79 -51 83 -37
rect 52 -55 83 -51
rect 52 -67 56 -55
rect 26 -71 56 -67
rect 26 -84 30 -71
<< labels >>
rlabel metal1 -30 20 -21 24 1 Vdd
rlabel space 122 -38 129 -33 1 Vdd
rlabel metal1 -30 -40 -23 -36 1 gnd
rlabel metal1 102 1 109 5 1 gnd
rlabel polycontact -23 -18 -19 -14 1 In_2
rlabel polycontact 45 42 49 46 1 In_2
rlabel pdcontact 18 27 22 47 1 In_2
rlabel ndcontact 18 -84 22 -74 1 In_2
rlabel polycontact 45 -54 49 -50 1 In_2
rlabel polycontact 19 14 23 18 1 In_1
rlabel polycontact 19 -71 23 -67 1 In_1
rlabel pdcontact 53 24 73 28 1 In_1
rlabel ndcontact 52 -47 62 -43 1 In_1
rlabel metal2 26 1 30 11 1 N1
rlabel metal2 26 27 30 47 1 N1
rlabel metal2 53 32 73 36 1 N1
rlabel metal2 26 -58 30 -38 1 N2
rlabel metal2 52 -55 62 -51 1 N2
rlabel metal2 26 -84 30 -74 1 N2
rlabel metal2 110 -37 114 -17 1 N2
rlabel metal2 103 13 107 17 1 N2
rlabel metal2 122 -14 126 -10 1 N1
rlabel metal2 118 1 122 11 1 N1
rlabel metal2 143 32 152 36 1 Out
rlabel metal2 -16 -31 -12 -21 1 N0
rlabel metal2 18 1 22 11 1 N0
rlabel metal2 -16 -5 -12 15 1 N0
rlabel metal2 18 -58 22 -38 1 N0
<< end >>
