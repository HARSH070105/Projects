magic
tech scmos
timestamp 1732055616
<< nwell >>
rect 0 0 24 34
<< ntransistor >>
rect 11 -19 13 -9
<< ptransistor >>
rect 11 6 13 26
<< ndiffusion >>
rect 10 -19 11 -9
rect 13 -19 14 -9
<< pdiffusion >>
rect 10 6 11 26
rect 13 6 14 26
<< ndcontact >>
rect 6 -19 10 -9
rect 14 -19 18 -9
<< pdcontact >>
rect 6 6 10 26
rect 14 6 18 26
<< polysilicon >>
rect 11 26 13 29
rect 11 -9 13 6
rect 11 -22 13 -19
<< polycontact >>
rect 7 -5 11 -1
<< metal1 >>
rect 0 34 24 38
rect 6 26 10 34
rect 14 -1 18 6
rect 0 -5 7 -1
rect 14 -5 24 -1
rect 14 -9 18 -5
rect 6 -23 10 -19
rect 0 -27 24 -23
<< labels >>
rlabel metal1 0 34 4 38 4 vdd
rlabel metal1 0 -5 4 -1 3 in
rlabel metal1 20 -5 24 -1 7 out
rlabel metal1 0 -27 4 -23 2 gnd
<< end >>
