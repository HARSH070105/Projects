* SPICE3 file created from xor1.ext - technology: scmos

.option scale=0.09u

M1000 a_25_n84# In_1 In_2 Gnd nfet w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M1001 a_53_31# In_2 In_1 w_45_18# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1002 a_25_1# In_1 a_18_1# Gnd nfet w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M1003 a_117_n37# a_115_n40# a_110_n37# w_104_n43# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1004 a_117_1# a_103_13# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=100 ps=60
M1005 a_25_n58# In_1 a_18_n58# w_12_n66# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1006 a_25_27# In_1 In_2 w_12_19# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1007 a_n17_n31# In_2 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1008 a_n17_n5# In_2 Vdd w_n30_n13# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1009 In_1 In_2 a_52_n55# Gnd nfet w=10 l=2
+  ad=50 pd=30 as=50 ps=30
C0 w_n30_n13# In_2 0.08fF
C1 w_12_19# In_1 0.08fF
C2 a_115_n40# N1 0.03fF
C3 a_18_1# N0 0.04fF
C4 In_2 N2 0.09fF
C5 a_25_27# N1 0.05fF
C6 w_12_n66# N2 0.21fF
C7 gnd a_n17_n31# 0.14fF
C8 In_2 a_52_n55# 0.05fF
C9 w_104_n43# N1 0.06fF
C10 a_117_1# gnd 0.10fF
C11 w_12_19# N1 0.21fF
C12 w_104_n43# a_110_n37# 0.03fF
C13 In_2 gnd 0.05fF
C14 w_104_n43# a_115_n40# 0.15fF
C15 In_1 In_2 0.08fF
C16 w_n30_n13# a_n17_n5# 0.03fF
C17 a_52_n55# N2 0.06fF
C18 w_12_19# a_25_27# 0.03fF
C19 w_12_n66# In_1 0.08fF
C20 w_45_18# In_2 0.13fF
C21 a_18_n58# N0 0.05fF
C22 a_n17_n31# N0 0.04fF
C23 a_18_n58# a_25_n58# 0.21fF
C24 a_117_1# N1 0.04fF
C25 a_143_32# N1 0.05fF
C26 a_103_13# N2 0.03fF
C27 In_2 N1 0.01fF
C28 w_12_n66# N0 0.19fF
C29 In_1 a_52_n55# 0.10fF
C30 w_n30_n13# N0 0.21fF
C31 w_12_n66# a_25_n58# 0.03fF
C32 In_1 gnd 0.03fF
C33 N0 N2 0.05fF
C34 In_1 a_25_1# 0.03fF
C35 In_1 a_53_31# 0.21fF
C36 In_2 a_25_27# 0.24fF
C37 w_n30_n13# Vdd 0.07fF
C38 w_45_18# a_53_31# 0.03fF
C39 a_25_n58# N2 0.05fF
C40 w_45_18# In_1 0.06fF
C41 w_12_19# In_2 0.07fF
C42 a_110_n37# N2 0.05fF
C43 a_n17_n5# N0 0.05fF
C44 a_110_n37# a_117_n37# 0.21fF
C45 a_25_1# N1 0.04fF
C46 a_53_31# N1 0.07fF
C47 w_104_n43# N2 0.19fF
C48 In_1 N0 0.26fF
C49 In_2 a_25_n84# 0.14fF
C50 w_45_18# N1 0.21fF
C51 Vdd a_n17_n5# 0.24fF
C52 w_12_n66# a_18_n58# 0.03fF
C53 w_104_n43# a_117_n37# 0.04fF
C54 a_18_1# a_25_1# 0.10fF
C55 In_1 a_18_1# 0.08fF
C56 N1 N0 0.03fF
C57 a_25_n84# N2 0.04fF
C58 N2 Gnd 0.54fF **FLOATING
C59 N0 Gnd 0.71fF **FLOATING
C60 a_25_n84# Gnd 0.02fF
C61 a_52_n55# Gnd 0.01fF
C62 a_117_n37# Gnd 0.01fF
C63 a_n17_n31# Gnd 0.02fF
C64 gnd Gnd 0.11fF
C65 a_103_13# Gnd 0.14fF
C66 a_143_32# Gnd 0.11fF **FLOATING
C67 In_2 Gnd 0.14fF
C68 In_1 Gnd 0.74fF
C69 w_104_n43# Gnd 0.82fF
C70 w_12_n66# Gnd 0.82fF
C71 w_45_18# Gnd 0.29fF
C72 w_12_19# Gnd 0.67fF
C73 w_n30_n13# Gnd 0.48fF
