magic
tech scmos
timestamp 1732101596
<< nwell >>
rect -6 19 18 131
<< ntransistor >>
rect 5 0 7 10
rect 21 0 23 10
<< ptransistor >>
rect 5 83 7 123
rect 5 25 7 65
<< ndiffusion >>
rect 4 0 5 10
rect 7 0 8 10
rect 20 0 21 10
rect 23 0 24 10
<< pdiffusion >>
rect 4 83 5 123
rect 7 83 8 123
rect 4 25 5 65
rect 7 25 8 65
<< ndcontact >>
rect 0 0 4 10
rect 8 0 12 10
rect 16 0 20 10
rect 24 0 28 10
<< pdcontact >>
rect 0 83 4 123
rect 8 83 12 123
rect 0 25 4 65
rect 8 25 12 65
<< polysilicon >>
rect 5 123 7 126
rect 5 76 7 83
rect 5 65 7 72
rect 5 22 7 25
rect 5 10 7 13
rect 21 10 23 28
rect 5 -7 7 0
rect 21 -3 23 0
<< polycontact >>
rect 1 76 5 80
rect 1 68 5 72
rect 23 24 27 28
rect 1 -7 5 -3
<< metal1 >>
rect -6 131 18 135
rect 0 123 4 131
rect -14 76 1 80
rect -14 -3 -11 76
rect 8 65 12 83
rect 0 18 4 25
rect 0 14 28 18
rect 0 10 4 14
rect 16 10 20 14
rect -14 -7 1 -3
rect 8 -10 12 0
rect 24 -10 28 0
rect -7 -14 28 -10
<< m2contact >>
rect -4 68 1 73
rect 23 28 28 33
<< metal2 >>
rect -10 68 -4 72
rect 1 68 27 72
rect 23 33 27 68
rect 23 24 27 28
<< labels >>
rlabel metal1 -6 -13 -4 -11 1 gnd
rlabel metal1 -5 132 -3 134 5 vdd
rlabel metal2 -9 69 -7 71 1 in2
rlabel metal1 25 15 27 17 7 out
rlabel metal1 -10 77 -8 79 3 in1
<< end >>
